** ICARIS generated Circuit **
r1 1 0 1
v2 1 0 dc 5
.END